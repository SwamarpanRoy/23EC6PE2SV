//------------------------------------------------------------------------------
//File       : dummy_dut.sv
//Author     : Swamarpan Roy/1BM23C305
//Created    : 2026-01-29
//Module     : dummy_dut
//Project    : SystemVerilog and Verification (23EC6PE2SV)
//Faculty    : Prof. Ajaykumar Devarapalli
//Description: A placeholder dummy DUT for the class-based Packet verification lab.
//------------------------------------------------------------------------------

module dummy_dut;
endmodule
